LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY JMP_DETECT_UNIT IS
	PORT (
		disable : IN STD_LOGIC;
		FLAGS_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		OT_CODE : IN STD_LOGIC_VECTOR(1 DOWNTO 0); --(OPERATIONAL TYPE)
		ID_CODE : IN STD_LOGIC_VECTOR(2 DOWNTO 0); --(Instruction identification)

		CHECK_JMP : OUT STD_LOGIC;
		FLAGS_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY JMP_DETECT_UNIT;
ARCHITECTURE ARCH_JMP_DETECT_UNIT OF JMP_DETECT_UNIT IS

	SIGNAL N_flag : STD_LOGIC; --(NEGATIVE FLAG)
	SIGNAL C_FLAG : STD_LOGIC; --(CARRAY FLAG)
	SIGNAL Z_flag : STD_LOGIC; --(ZERO FLAG)
BEGIN

	-- HERE WE CHECK IF THIS IS A JUMP INSTRUCTION
	CHECK_JMP <= '1' WHEN ((OT_CODE = "11") AND (ID_CODE = "100"))
		ELSE
		'1' WHEN ((OT_CODE = "11") AND (ID_CODE = "000") AND (FLAGS_IN(0) = '1'))
		ELSE
		'1' WHEN ((OT_CODE = "11") AND (ID_CODE = "001") AND (FLAGS_IN(2) = '1'))
		ELSE
		'1' WHEN ((OT_CODE = "11") AND (ID_CODE = "010") AND (FLAGS_IN(1) = '1'))
		ELSE
		'1' WHEN ((OT_CODE = "11") AND (ID_CODE = "011"))
		ELSE
		'0' WHEN disable = '1'
		ELSE
		'0';

	--ZERO JUMP INSTRUCTION
	Z_flag <= '0' WHEN ((OT_CODE = "11") AND (ID_CODE = "000") AND (FLAGS_IN(0) = '1'))
		ELSE
		FLAGS_IN(0);

	--NEGATIVE JUMP INSTRUCTION
	N_flag <= '0' WHEN ((OT_CODE = "11") AND (ID_CODE = "001") AND (FLAGS_IN(1) = '1'))
		ELSE
		FLAGS_IN(1);

	--CARRY JUMP INSTRUCTION
	C_FLAG <= '0' WHEN ((OT_CODE = "11") AND (ID_CODE = "010") AND (FLAGS_IN(2) = '1'))
		ELSE
		FLAGS_IN(2);
	FLAGS_OUT <= '0' & C_FLAG & N_flag & Z_flag;

END ARCH_JMP_DETECT_UNIT;